always_ff @( clock ) begin : blockName
    case
        
    endcase
end
always_comb begin : tea
    a = 
end
// a is a variable
reg k; // after comment

always_comb begin
    k = 33;
end

toInst u_toInst(
	.a(a),
    .b(b),
    .c(c)
);

toInst 
#(
    .width(width),
    .width2(width2)
)
u_toInst(
	.a(a),
    .b(b),
    .c(c)
);

mod_name instance_name (.*);
toInst 
#(
    .width_sdajdads (width_sdajdads ),
    .width2_asdf    (width2_asdf    )
)
u_toInst(
	.aasdasd     (aasdasd     ),
    .bdasdasf    (bdasdasf    ),
    .cfafafafasf (cfafafafasf )
);

/*
dasdas
dasda
*/
// sdas
  reg aa  = 15; 
  reg aaa = 33; 

  wire   [13:fd 0] aa          ;      
  wire   [13:   0] bb          ;      
  wire   [13:   0] vv          ;      
  reg    [12:   0] dd  [35:15] ;      
  assign a = 15    
  assign b = 35848 


always_comb begin
  a      = 15     ; 
  addfdf = 33     ; 
  fff    = 15+gfdg; 
end

always_ff(@posedge clk)begin
  a    <= 57; 
  c    <= df; 
  fsdf <= df; 
    if(fsdfsd)begin
        dfdsf <= df; 
    end
    else begin
        dfsdf <=fdfdsfsfs;
        fdsfds <= dsfsdfs;
    end
end

aa
toInst 
#(
    .width_sdajdads (width_sdajdads ),
    .width2_asdf    (width2_asdf    )
)
u_toInst(
	.aasdasd     (aasdasd     ),
    .bdasdasf    (bdasdasf    ),
    .cfafafafasf (cfafafafasf )
);

